
module cpu 
(
);




endmodule
